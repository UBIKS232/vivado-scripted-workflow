module top();

endmodule

