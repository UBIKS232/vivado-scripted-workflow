module tb_test();

endmodule
