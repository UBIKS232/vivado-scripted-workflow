1ns/1ps
module tb_test();

endmodule
