`timescale 1ns / 1ps

module tb_top();

	/*iverilog */
	initial
	begin
		("tb_top.vcd");
		(0, tb_top);
	end
	/*iverilog */


endmodule

